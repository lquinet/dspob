PLL_BUF_inst : PLL_BUF PORT MAP (
		areset	 => areset_sig,
		inclk0	 => inclk0_sig,
		c0	 => c0_sig
	);
